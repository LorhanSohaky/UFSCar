library verilog;
use verilog.vl_types.all;
entity decodificador_TB is
end decodificador_TB;
