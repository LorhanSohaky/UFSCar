library verilog;
use verilog.vl_types.all;
entity Etapa1_vlg_vec_tst is
end Etapa1_vlg_vec_tst;
