library verilog;
use verilog.vl_types.all;
entity separa is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        E               : in     vl_logic;
        z0              : out    vl_logic;
        z1              : out    vl_logic;
        z2              : out    vl_logic;
        z3              : out    vl_logic;
        z4              : out    vl_logic
    );
end separa;
