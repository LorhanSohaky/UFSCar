module regn ( R, Rin, Clock, Q );
  parameter n = 8;

  input [n-1:0] R;
  input Rin, Clock;

  output [n-1:0] Q;
  reg [n-1:0] Q;

  always @( posedge Clock )
    if ( Rin )
      Q <= R;
endmodule
