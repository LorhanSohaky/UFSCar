library verilog;
use verilog.vl_types.all;
entity MeioSomador4Bits_vlg_vec_tst is
end MeioSomador4Bits_vlg_vec_tst;
