library verilog;
use verilog.vl_types.all;
entity maquina_TB is
end maquina_TB;
