library verilog;
use verilog.vl_types.all;
entity circuitoAdicional_TB is
end circuitoAdicional_TB;
