library verilog;
use verilog.vl_types.all;
entity Projeto2_vlg_check_tst is
    port(
        LEDG            : in     vl_logic_vector(1 downto 1);
        sampler_rx      : in     vl_logic
    );
end Projeto2_vlg_check_tst;
