library verilog;
use verilog.vl_types.all;
entity Etapa2_vlg_vec_tst is
end Etapa2_vlg_vec_tst;
