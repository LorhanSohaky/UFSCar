library verilog;
use verilog.vl_types.all;
entity projetoPessoal_TB is
end projetoPessoal_TB;
