library verilog;
use verilog.vl_types.all;
entity tcounter is
end tcounter;
