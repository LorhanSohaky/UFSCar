library verilog;
use verilog.vl_types.all;
entity Projeto2_vlg_vec_tst is
end Projeto2_vlg_vec_tst;
